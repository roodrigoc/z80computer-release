

localparam [16383:0] fontmem_new = {
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00111100,
8'b00111100,
8'b00111100,
8'b00111100,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00011110,
8'b00000110,
8'b00001100,
8'b00011000,
8'b00001110,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110110,
8'b00110110,
8'b00110110,
8'b00011110,

8'b00111000,
8'b00111100,
8'b00110110,
8'b00110111,
8'b00110000,
8'b00110000,
8'b00110000,
8'b11110000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00011000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00011000,
8'b00011000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00011100,
8'b00110110,
8'b00110110,
8'b00011100,

8'b00000000,
8'b00000000,
8'b00111011,
8'b01101110,
8'b00000000,
8'b00111011,
8'b01101110,
8'b00000000,

8'b00000000,
8'b00001100,
8'b00001100,
8'b00000000,
8'b00111111,
8'b00000000,
8'b00001100,
8'b00001100,

8'b00001110,
8'b00011011,
8'b00011011,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,

8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b11011000,
8'b11011000,
8'b01110000,

8'b00000000,
8'b00111111,
8'b00000000,
8'b00011000,
8'b00001100,
8'b00000110,
8'b00001100,
8'b00011000,

8'b00000000,
8'b00111111,
8'b00000000,
8'b00000110,
8'b00001100,
8'b00011000,
8'b00001100,
8'b00000110,

8'b00000000,
8'b00111111,
8'b00000000,
8'b00001100,
8'b00001100,
8'b00111111,
8'b00001100,
8'b00001100,

8'b00000000,
8'b00000000,
8'b00111111,
8'b00000000,
8'b00111111,
8'b00000000,
8'b00111111,
8'b00000000,

8'b00000000,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00011110,

8'b00000000,
8'b00011100,
8'b00000110,
8'b00000011,
8'b00011111,
8'b00000011,
8'b00000110,
8'b00011100,

8'b00000011,
8'b00000110,
8'b01111110,
8'b11011011,
8'b11011011,
8'b01111110,
8'b00110000,
8'b01100000,

8'b00000000,
8'b00000000,
8'b01111110,
8'b11011011,
8'b11011011,
8'b01111110,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00111110,
8'b00011000,
8'b00001100,
8'b00111000,

8'b00000000,
8'b01110111,
8'b00110110,
8'b00110110,
8'b01100011,
8'b01100011,
8'b00110110,
8'b00011100,

8'b00000000,
8'b00011100,
8'b00110110,
8'b01100011,
8'b01111111,
8'b01100011,
8'b00110110,
8'b00011100,

8'b00111111,
8'b00001100,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00011110,
8'b00001100,
8'b00111111,

8'b00000000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00111011,
8'b01101110,
8'b00000000,

8'b00000011,
8'b00000110,
8'b00111110,
8'b01100110,
8'b01100110,
8'b01100110,
8'b01100110,
8'b00000000,

8'b00000000,
8'b00001110,
8'b00011011,
8'b00011011,
8'b00011011,
8'b01111110,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00111111,
8'b00110011,
8'b00000110,
8'b00001100,
8'b00000110,
8'b00110011,
8'b00111111,

8'b00000000,
8'b00110110,
8'b00110110,
8'b00110110,
8'b00110110,
8'b00110110,
8'b01111111,
8'b00000000,

8'b00000000,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00110011,
8'b00111111,
8'b00000000,

8'b00000011,
8'b00000011,
8'b00011111,
8'b00110011,
8'b00011111,
8'b00110011,
8'b00011110,
8'b00000000,

8'b00000000,
8'b01101110,
8'b00111011,
8'b00010011,
8'b00111011,
8'b01101110,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,

8'b11110000,
8'b11110000,
8'b11110000,
8'b11110000,
8'b11110000,
8'b11110000,
8'b11110000,
8'b11110000,

8'b00001111,
8'b00001111,
8'b00001111,
8'b00001111,
8'b00001111,
8'b00001111,
8'b00001111,
8'b00001111,

8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,

8'b00011000,
8'b00011000,
8'b00011000,
8'b11111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00011111,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,

8'b00011000,
8'b00011000,
8'b00011000,
8'b11111111,
8'b00011000,
8'b11111111,
8'b00011000,
8'b00011000,

8'b01101100,
8'b01101100,
8'b01101100,
8'b11111111,
8'b01101100,
8'b01101100,
8'b01101100,
8'b01101100,

8'b01101100,
8'b01101100,
8'b01101100,
8'b11111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00011000,
8'b00011000,
8'b00011000,
8'b11111000,
8'b00011000,
8'b11111000,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b11111000,
8'b00011000,
8'b11111000,
8'b00011000,
8'b00011000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b11111100,
8'b01101100,
8'b01101100,
8'b01101100,
8'b01101100,

8'b01101100,
8'b01101100,
8'b01101100,
8'b11111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00011000,
8'b00011000,
8'b00011000,
8'b11111111,
8'b00000000,
8'b11111111,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b11111111,
8'b01101100,
8'b01101100,
8'b01101100,
8'b01101100,

8'b00000000,
8'b00000000,
8'b00000000,
8'b11111111,
8'b00000000,
8'b11111111,
8'b00011000,
8'b00011000,

8'b01101100,
8'b01101100,
8'b01101100,
8'b11101111,
8'b00000000,
8'b11101111,
8'b01101100,
8'b01101100,

8'b00000000,
8'b00000000,
8'b00000000,
8'b11111111,
8'b00000000,
8'b11111111,
8'b00000000,
8'b00000000,

8'b01101100,
8'b01101100,
8'b01101100,
8'b11101100,
8'b00001100,
8'b11101100,
8'b01101100,
8'b01101100,

8'b01101100,
8'b01101100,
8'b01101100,
8'b11101111,
8'b00000000,
8'b11111111,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b11111111,
8'b00000000,
8'b11101111,
8'b01101100,
8'b01101100,

8'b01101100,
8'b01101100,
8'b01101100,
8'b11101100,
8'b00001100,
8'b11111100,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b11111100,
8'b00001100,
8'b11101100,
8'b01101100,
8'b01101100,

8'b01101100,
8'b01101100,
8'b01101100,
8'b11101100,
8'b01101100,
8'b01101100,
8'b01101100,
8'b01101100,

8'b00011000,
8'b00011000,
8'b00011000,
8'b11111000,
8'b00011000,
8'b11111000,
8'b00011000,
8'b00011000,

8'b00011000,
8'b00011000,
8'b00011000,
8'b11111111,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b11111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00011000,
8'b00011000,
8'b00011000,
8'b11111000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,

8'b00011000,
8'b00011000,
8'b00011000,
8'b11111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b11111111,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b11111000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,

8'b00011000,
8'b00011000,
8'b00011000,
8'b00011111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00011111,
8'b00011000,
8'b00011111,
8'b00011000,
8'b00011000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b01111111,
8'b01101100,
8'b01101100,
8'b01101100,
8'b01101100,

8'b00000000,
8'b00000000,
8'b00000000,
8'b01111111,
8'b01100000,
8'b01101111,
8'b01101100,
8'b01101100,

8'b01101100,
8'b01101100,
8'b01101100,
8'b01101111,
8'b01100000,
8'b01111111,
8'b00000000,
8'b00000000,

8'b01101100,
8'b01101100,
8'b01101100,
8'b01101100,
8'b01101100,
8'b01101100,
8'b01101100,
8'b01101100,

8'b01101100,
8'b01101100,
8'b01101100,
8'b01101111,
8'b01100000,
8'b01101111,
8'b01101100,
8'b01101100,

8'b00011000,
8'b00011000,
8'b00011000,
8'b00011111,
8'b00011000,
8'b00011111,
8'b00000000,
8'b00000000,

8'b01101100,
8'b01101100,
8'b01101100,
8'b01111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b01101100,
8'b01101100,
8'b01101100,
8'b01101111,
8'b01101100,
8'b01101100,
8'b01101100,
8'b01101100,

8'b00011000,
8'b00011000,
8'b00011000,
8'b00011111,
8'b00011000,
8'b00011111,
8'b00011000,
8'b00011000,

8'b00011000,
8'b00011000,
8'b00011000,
8'b00011111,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,

8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,

8'b01110111,
8'b11011011,
8'b11101110,
8'b11011011,
8'b01110111,
8'b11011011,
8'b11101110,
8'b11011011,

8'b01010101,
8'b10101010,
8'b01010101,
8'b10101010,
8'b01010101,
8'b10101010,
8'b01010101,
8'b10101010,

8'b00010001,
8'b01000100,
8'b00010001,
8'b01000100,
8'b00010001,
8'b01000100,
8'b00010001,
8'b01000100,

8'b00000000,
8'b00000000,
8'b00110011,
8'b01100110,
8'b11001100,
8'b01100110,
8'b00110011,
8'b00000000,

8'b00000000,
8'b00000000,
8'b11001100,
8'b01100110,
8'b00110011,
8'b01100110,
8'b11001100,
8'b00000000,

8'b00000000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00000000,
8'b00011000,
8'b00011000,

8'b11000000,
8'b11110011,
8'b11110110,
8'b11101100,
8'b11011011,
8'b00110011,
8'b01100011,
8'b11000011,

8'b11110000,
8'b00110011,
8'b01100110,
8'b11001100,
8'b01111011,
8'b00110011,
8'b01100011,
8'b11000011,

8'b00000000,
8'b00000000,
8'b00110000,
8'b00110000,
8'b00111111,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000011,
8'b00000011,
8'b00111111,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00000011,
8'b00000110,
8'b00001100,
8'b00000000,
8'b00001100,

8'b00000000,
8'b00000000,
8'b00111110,
8'b00000000,
8'b00011100,
8'b00110110,
8'b00110110,
8'b00011100,

8'b00000000,
8'b00000000,
8'b01111110,
8'b00000000,
8'b01111100,
8'b00110110,
8'b00110110,
8'b00111100,

8'b00000000,
8'b00110011,
8'b00111011,
8'b00111111,
8'b00110111,
8'b00110011,
8'b00000000,
8'b00111111,

8'b00000000,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00011111,
8'b00000000,
8'b00011111,
8'b00000000,

8'b00000000,
8'b01111110,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00000000,
8'b00111000,
8'b00000000,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00011110,
8'b00000000,
8'b00111000,
8'b00000000,

8'b00000000,
8'b00011110,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001110,
8'b00000000,
8'b00011100,

8'b00000000,
8'b01111110,
8'b00110011,
8'b00111110,
8'b00110000,
8'b00011110,
8'b00000000,
8'b00111000,

8'b00001110,
8'b00011011,
8'b00011000,
8'b00011000,
8'b00111100,
8'b00011000,
8'b11011000,
8'b01110000,

8'b11100011,
8'b01100011,
8'b11110011,
8'b01100011,
8'b01011111,
8'b00110011,
8'b00110011,
8'b00011111,

8'b00001100,
8'b00001100,
8'b00111111,
8'b00001100,
8'b00111111,
8'b00011110,
8'b00110011,
8'b00110011,

8'b00000000,
8'b00111111,
8'b01100111,
8'b00000110,
8'b00001111,
8'b00100110,
8'b00110110,
8'b00011100,

8'b00011000,
8'b00011000,
8'b01111110,
8'b00000011,
8'b00000011,
8'b01111110,
8'b00011000,
8'b00011000,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00000000,
8'b00110011,

8'b00000000,
8'b00011000,
8'b00111100,
8'b01100110,
8'b01100110,
8'b00111100,
8'b00011000,
8'b11000011,

8'b00011111,
8'b00110000,
8'b00111110,
8'b00110011,
8'b00110011,
8'b00000000,
8'b00110011,
8'b00000000,

8'b00000000,
8'b01111110,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00000000,
8'b00000111,
8'b00000000,

8'b00000000,
8'b01111110,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00000000,
8'b00110011,
8'b00011110,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00011110,
8'b00000000,
8'b00000111,
8'b00000000,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00011110,
8'b00000000,
8'b00110011,
8'b00000000,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00011110,
8'b00000000,
8'b00110011,
8'b00011110,

8'b00000000,
8'b01110011,
8'b00110011,
8'b00110011,
8'b01111111,
8'b00110011,
8'b00110110,
8'b01111100,

8'b00000000,
8'b11111110,
8'b00110011,
8'b11111110,
8'b00110000,
8'b11111110,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00111111,
8'b00000110,
8'b00011110,
8'b00000110,
8'b00111111,
8'b00000000,
8'b00111000,

8'b00000000,
8'b00110011,
8'b00111111,
8'b00110011,
8'b00011110,
8'b00000000,
8'b00001100,
8'b00001100,

8'b00000000,
8'b01100011,
8'b01100011,
8'b01111111,
8'b01100011,
8'b00110110,
8'b00011100,
8'b01100011,

8'b00000000,
8'b00011110,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001110,
8'b00000000,
8'b00000111,

8'b00000000,
8'b00111100,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011100,
8'b01100011,
8'b00111110,

8'b00000000,
8'b00011110,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001110,
8'b00000000,
8'b00110011,

8'b00000000,
8'b00011110,
8'b00000011,
8'b00111111,
8'b00110011,
8'b00011110,
8'b00000000,
8'b00000111,

8'b00000000,
8'b00011110,
8'b00000011,
8'b00111111,
8'b00110011,
8'b00011110,
8'b00000000,
8'b00110011,

8'b00000000,
8'b00111100,
8'b00000110,
8'b01111110,
8'b01100110,
8'b00111100,
8'b11000011,
8'b01111110,

8'b00011100,
8'b00110000,
8'b00011110,
8'b00000011,
8'b00000011,
8'b00011110,
8'b00000000,
8'b00000000,

8'b00000000,
8'b01111110,
8'b00110011,
8'b00111110,
8'b00110000,
8'b00011110,
8'b00001100,
8'b00001100,

8'b00000000,
8'b01111110,
8'b00110011,
8'b00111110,
8'b00110000,
8'b00011110,
8'b00000000,
8'b00000111,

8'b00000000,
8'b01111110,
8'b00110011,
8'b00111110,
8'b00110000,
8'b00011110,
8'b00000000,
8'b00110011,

8'b00000000,
8'b11111100,
8'b01100110,
8'b01111100,
8'b01100000,
8'b00111100,
8'b11000011,
8'b01111110,

8'b00000000,
8'b00011110,
8'b00000011,
8'b00111111,
8'b00110011,
8'b00011110,
8'b00000000,
8'b00111000,

8'b00000000,
8'b01111110,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00000000,
8'b00110011,
8'b00000000,

8'b00011110,
8'b00110000,
8'b00011000,
8'b00011110,
8'b00110011,
8'b00000011,
8'b00110011,
8'b00011110,

8'b00000000,
8'b01111111,
8'b01100011,
8'b01100011,
8'b00110110,
8'b00011100,
8'b00001000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111011,
8'b01101110,

8'b00000000,
8'b00000111,
8'b00001100,
8'b00001100,
8'b00111000,
8'b00001100,
8'b00001100,
8'b00000111,

8'b00000000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00000000,
8'b00011000,
8'b00011000,
8'b00011000,

8'b00000000,
8'b00111000,
8'b00001100,
8'b00001100,
8'b00000111,
8'b00001100,
8'b00001100,
8'b00111000,

8'b00000000,
8'b00111111,
8'b00100110,
8'b00001100,
8'b00011001,
8'b00111111,
8'b00000000,
8'b00000000,

8'b00011111,
8'b00110000,
8'b00111110,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00000000,
8'b00000000,

8'b00000000,
8'b01100011,
8'b00110110,
8'b00011100,
8'b00110110,
8'b01100011,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00110110,
8'b01111111,
8'b01111111,
8'b01101011,
8'b01100011,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00001100,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00000000,
8'b00000000,

8'b00000000,
8'b01101110,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00011000,
8'b00101100,
8'b00001100,
8'b00001100,
8'b00111110,
8'b00001100,
8'b00001000,

8'b00000000,
8'b00011111,
8'b00110000,
8'b00011110,
8'b00000011,
8'b00111110,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00001111,
8'b00000110,
8'b01100110,
8'b01101110,
8'b00111011,
8'b00000000,
8'b00000000,

8'b01111000,
8'b00110000,
8'b00111110,
8'b00110011,
8'b00110011,
8'b01101110,
8'b00000000,
8'b00000000,

8'b00001111,
8'b00000110,
8'b00111110,
8'b01100110,
8'b01100110,
8'b00111011,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00011110,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00011111,
8'b00000000,
8'b00000000,

8'b00000000,
8'b01100011,
8'b01101011,
8'b01111111,
8'b01111111,
8'b00110011,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00011110,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001110,

8'b00000000,
8'b01100111,
8'b00110110,
8'b00011110,
8'b00110110,
8'b01100110,
8'b00000110,
8'b00000111,

8'b00011110,
8'b00110011,
8'b00110011,
8'b00110000,
8'b00110000,
8'b00110000,
8'b00000000,
8'b00110000,

8'b00000000,
8'b00011110,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001110,
8'b00000000,
8'b00001100,

8'b00000000,
8'b01100111,
8'b01100110,
8'b01100110,
8'b01101110,
8'b00110110,
8'b00000110,
8'b00000111,

8'b00011111,
8'b00110000,
8'b00111110,
8'b00110011,
8'b00110011,
8'b01101110,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00001111,
8'b00000110,
8'b00000110,
8'b00001111,
8'b00000110,
8'b00110110,
8'b00011100,

8'b00000000,
8'b00011110,
8'b00000011,
8'b00111111,
8'b00110011,
8'b00011110,
8'b00000000,
8'b00000000,

8'b00000000,
8'b01101110,
8'b00110011,
8'b00110011,
8'b00111110,
8'b00110000,
8'b00110000,
8'b00111000,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00000011,
8'b00110011,
8'b00011110,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00111011,
8'b01100110,
8'b01100110,
8'b00111110,
8'b00000110,
8'b00000110,
8'b00000111,

8'b00000000,
8'b01101110,
8'b00110011,
8'b00111110,
8'b00110000,
8'b00011110,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00011000,
8'b00001100,
8'b00001100,

8'b11111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01100011,
8'b00110110,
8'b00011100,
8'b00001000,

8'b00000000,
8'b00011110,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011110,

8'b00000000,
8'b01000000,
8'b01100000,
8'b00110000,
8'b00011000,
8'b00001100,
8'b00000110,
8'b00000011,

8'b00000000,
8'b00011110,
8'b00000110,
8'b00000110,
8'b00000110,
8'b00000110,
8'b00000110,
8'b00011110,

8'b00000000,
8'b01111111,
8'b01100110,
8'b01001100,
8'b00011000,
8'b00110001,
8'b01100011,
8'b01111111,

8'b00000000,
8'b00011110,
8'b00001100,
8'b00001100,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00110011,

8'b00000000,
8'b01100011,
8'b00110110,
8'b00011100,
8'b00011100,
8'b00110110,
8'b01100011,
8'b01100011,

8'b00000000,
8'b01100011,
8'b01110111,
8'b01111111,
8'b01101011,
8'b01100011,
8'b01100011,
8'b01100011,

8'b00000000,
8'b00001100,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00110011,

8'b00000000,
8'b00111111,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00110011,

8'b00000000,
8'b00011110,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00101101,
8'b00111111,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00111000,
8'b00001110,
8'b00000111,
8'b00110011,
8'b00011110,

8'b00000000,
8'b01100111,
8'b01100110,
8'b00110110,
8'b00111110,
8'b01100110,
8'b01100110,
8'b00111111,

8'b00000000,
8'b00111000,
8'b00011110,
8'b00111011,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00011110,

8'b00000000,
8'b00001111,
8'b00000110,
8'b00000110,
8'b00111110,
8'b01100110,
8'b01100110,
8'b00111111,

8'b00000000,
8'b00011100,
8'b00110110,
8'b01100011,
8'b01100011,
8'b01100011,
8'b00110110,
8'b00011100,

8'b00000000,
8'b01100011,
8'b01100011,
8'b01110011,
8'b01111011,
8'b01101111,
8'b01100111,
8'b01100011,

8'b00000000,
8'b01100011,
8'b01100011,
8'b01101011,
8'b01111111,
8'b01111111,
8'b01110111,
8'b01100011,

8'b00000000,
8'b01111111,
8'b01100110,
8'b01000110,
8'b00000110,
8'b00000110,
8'b00000110,
8'b00001111,

8'b00000000,
8'b01100111,
8'b01100110,
8'b00110110,
8'b00011110,
8'b00110110,
8'b01100110,
8'b01100111,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00110000,
8'b00110000,
8'b00110000,
8'b01111000,

8'b00000000,
8'b00011110,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00011110,

8'b00000000,
8'b00110011,
8'b00110011,
8'b00110011,
8'b00111111,
8'b00110011,
8'b00110011,
8'b00110011,

8'b00000000,
8'b01111100,
8'b01100110,
8'b01110011,
8'b00000011,
8'b00000011,
8'b01100110,
8'b00111100,

8'b00000000,
8'b00001111,
8'b00000110,
8'b00010110,
8'b00011110,
8'b00010110,
8'b01000110,
8'b01111111,

8'b00000000,
8'b01111111,
8'b01000110,
8'b00010110,
8'b00011110,
8'b00010110,
8'b01000110,
8'b01111111,

8'b00000000,
8'b00011111,
8'b00110110,
8'b01100110,
8'b01100110,
8'b01100110,
8'b00110110,
8'b00011111,

8'b00000000,
8'b00111100,
8'b01100110,
8'b00000011,
8'b00000011,
8'b00000011,
8'b01100110,
8'b00111100,

8'b00000000,
8'b00111111,
8'b01100110,
8'b01100110,
8'b00111110,
8'b01100110,
8'b01100110,
8'b00111111,

8'b00000000,
8'b00110011,
8'b00110011,
8'b00111111,
8'b00110011,
8'b00110011,
8'b00011110,
8'b00001100,

8'b00000000,
8'b00011110,
8'b00000011,
8'b01111011,
8'b01111011,
8'b01111011,
8'b01100011,
8'b00111110,

8'b00000000,
8'b00001100,
8'b00000000,
8'b00001100,
8'b00011000,
8'b00110000,
8'b00110011,
8'b00011110,

8'b00000000,
8'b00000110,
8'b00001100,
8'b00011000,
8'b00110000,
8'b00011000,
8'b00001100,
8'b00000110,

8'b00000000,
8'b00000000,
8'b00111111,
8'b00000000,
8'b00000000,
8'b00111111,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00011000,
8'b00001100,
8'b00000110,
8'b00000011,
8'b00000110,
8'b00001100,
8'b00011000,

8'b00000110,
8'b00001100,
8'b00001100,
8'b00000000,
8'b00000000,
8'b00001100,
8'b00001100,
8'b00000000,

8'b00000000,
8'b00001100,
8'b00001100,
8'b00000000,
8'b00000000,
8'b00001100,
8'b00001100,
8'b00000000,

8'b00000000,
8'b00001110,
8'b00011000,
8'b00110000,
8'b00111110,
8'b00110011,
8'b00110011,
8'b00011110,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00011110,

8'b00000000,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00011000,
8'b00110000,
8'b00110011,
8'b00111111,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00110011,
8'b00011111,
8'b00000011,
8'b00000110,
8'b00011100,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00110000,
8'b00110000,
8'b00011111,
8'b00000011,
8'b00111111,

8'b00000000,
8'b01111000,
8'b00110000,
8'b01111111,
8'b00110011,
8'b00110110,
8'b00111100,
8'b00111000,

8'b00000000,
8'b00011110,
8'b00110011,
8'b00110000,
8'b00011100,
8'b00110000,
8'b00110011,
8'b00011110,

8'b00000000,
8'b00111111,
8'b00110011,
8'b00000110,
8'b00011100,
8'b00110000,
8'b00110011,
8'b00011110,

8'b00000000,
8'b00111111,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001110,
8'b00001100,

8'b00000000,
8'b00111110,
8'b01100111,
8'b01101111,
8'b01111011,
8'b01110011,
8'b01100011,
8'b00111110,

8'b00000000,
8'b00000001,
8'b00000011,
8'b00000110,
8'b00001100,
8'b00011000,
8'b00110000,
8'b01100000,

8'b00000000,
8'b00001100,
8'b00001100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111111,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00000110,
8'b00001100,
8'b00001100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00001100,
8'b00001100,
8'b00111111,
8'b00001100,
8'b00001100,
8'b00000000,

8'b00000000,
8'b00000000,
8'b01100110,
8'b00111100,
8'b11111111,
8'b00111100,
8'b01100110,
8'b00000000,

8'b00000000,
8'b00000110,
8'b00001100,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00001100,
8'b00000110,

8'b00000000,
8'b00011000,
8'b00001100,
8'b00000110,
8'b00000110,
8'b00000110,
8'b00001100,
8'b00011000,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000110,
8'b00000110,

8'b00000000,
8'b01101110,
8'b00110011,
8'b00111011,
8'b01101110,
8'b00011100,
8'b00110110,
8'b00011100,

8'b00000000,
8'b01100011,
8'b01100110,
8'b00001100,
8'b00011000,
8'b00110011,
8'b01100011,
8'b00000000,

8'b00000000,
8'b00001100,
8'b00011111,
8'b00110000,
8'b00011110,
8'b00000011,
8'b00111110,
8'b00001100,

8'b00000000,
8'b00110110,
8'b00110110,
8'b01111111,
8'b00110110,
8'b01111111,
8'b00110110,
8'b00110110,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110110,
8'b00110110,

8'b00000000,
8'b00001100,
8'b00000000,
8'b00001100,
8'b00001100,
8'b00011110,
8'b00011110,
8'b00001100,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00011000,
8'b00111100,
8'b01111110,
8'b11111111,
8'b11111111,
8'b00000000,

8'b00000000,
8'b00000000,
8'b11111111,
8'b11111111,
8'b01111110,
8'b00111100,
8'b00011000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00100100,
8'b01100110,
8'b11111111,
8'b01100110,
8'b00100100,
8'b00000000,

8'b00000000,
8'b00000000,
8'b01111111,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00001100,
8'b00000110,
8'b01111111,
8'b00000110,
8'b00001100,
8'b00000000,

8'b00000000,
8'b00000000,
8'b00011000,
8'b00110000,
8'b01111111,
8'b00110000,
8'b00011000,
8'b00000000,

8'b00000000,
8'b00011000,
8'b00111100,
8'b01111110,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,

8'b00000000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b01111110,
8'b00111100,
8'b00011000,

8'b11111111,
8'b00011000,
8'b00111100,
8'b01111110,
8'b00011000,
8'b01111110,
8'b00111100,
8'b00011000,

8'b00000000,
8'b01111110,
8'b01111110,
8'b01111110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,

8'b00011110,
8'b00110011,
8'b00011100,
8'b00110110,
8'b00110110,
8'b00011100,
8'b11000110,
8'b01111100,

8'b00000000,
8'b11011000,
8'b11011000,
8'b11011000,
8'b11011110,
8'b11011011,
8'b11011011,
8'b11111110,

8'b00000000,
8'b01100110,
8'b00000000,
8'b01100110,
8'b01100110,
8'b01100110,
8'b01100110,
8'b01100110,

8'b00011000,
8'b00111100,
8'b01111110,
8'b00011000,
8'b00011000,
8'b01111110,
8'b00111100,
8'b00011000,

8'b00000000,
8'b01000000,
8'b01110000,
8'b01111100,
8'b01111111,
8'b01111100,
8'b01110000,
8'b01000000,

8'b00000000,
8'b00000001,
8'b00000111,
8'b00011111,
8'b01111111,
8'b00011111,
8'b00000111,
8'b00000001,

8'b10011001,
8'b01011010,
8'b00111100,
8'b11100111,
8'b11100111,
8'b00111100,
8'b01011010,
8'b10011001,

8'b00000011,
8'b01100111,
8'b11100110,
8'b11000110,
8'b11000110,
8'b11111110,
8'b11000110,
8'b11111110,

8'b00000111,
8'b00001111,
8'b00001110,
8'b00001100,
8'b00001100,
8'b11111100,
8'b11001100,
8'b11111100,

8'b00011000,
8'b01111110,
8'b00011000,
8'b00111100,
8'b01100110,
8'b01100110,
8'b01100110,
8'b00111100,

8'b00011110,
8'b00110011,
8'b00110011,
8'b00110011,
8'b10111110,
8'b11110000,
8'b11100000,
8'b11110000,

8'b11111111,
8'b11000011,
8'b10011001,
8'b10111101,
8'b10111101,
8'b10011001,
8'b11000011,
8'b11111111,

8'b00000000,
8'b00111100,
8'b01100110,
8'b01000010,
8'b01000010,
8'b01100110,
8'b00111100,
8'b00000000,

8'b11111111,
8'b11111111,
8'b11100111,
8'b11000011,
8'b11000011,
8'b11100111,
8'b11111111,
8'b11111111,

8'b00000000,
8'b00000000,
8'b00011000,
8'b00111100,
8'b00111100,
8'b00011000,
8'b00000000,
8'b00000000,

8'b00111110,
8'b00011100,
8'b00111110,
8'b01111111,
8'b00111110,
8'b00011100,
8'b00001000,
8'b00001000,

8'b00111110,
8'b00011100,
8'b00111110,
8'b01111111,
8'b01111111,
8'b00011100,
8'b00111110,
8'b00011100,

8'b00000000,
8'b00001000,
8'b00011100,
8'b00111110,
8'b01111111,
8'b00111110,
8'b00011100,
8'b00001000,

8'b00000000,
8'b00001000,
8'b00011100,
8'b00111110,
8'b01111111,
8'b01111111,
8'b01111111,
8'b00110110,

8'b01111110,
8'b11111111,
8'b11100111,
8'b11000011,
8'b11111111,
8'b11011011,
8'b11111111,
8'b01111110,

8'b01111110,
8'b10000001,
8'b10011001,
8'b10111101,
8'b10000001,
8'b10100101,
8'b10000001,
8'b01111110,

8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000
};
